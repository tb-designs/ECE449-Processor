library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity PCincr is 
  port();

end PCincr;

architecture Behavioral of PCincr is


  end Behavioral;