----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 02/24/2020 04:18:32 PM
-- Design Name: 
-- Module Name: datapath - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library ieee;
use ieee.std_logic_1164.all;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
use ieee.numeric_std.all;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity processor is
    port ( --Inputs
        clk : in std_logic;
        sw_in : in std_logic_vector(1 downto 0);
        an_out : out std_logic_vector(3 downto 0);
        sseg_out : out std_logic_vector(6 downto 0);
        in_port : in std_logic_vector(9 downto 0);
        out_port : out std_logic
    );
end processor;

architecture behavioral of processor is

--Program Counter
component pc is
    port (
        clk : in std_logic;
        rst : in std_logic;
        pc_in : in std_logic_vector(15 downto 0);
        pc_out : out std_logic_vector(15 downto 0)  
    );
end component;

-- Memory Interface
component mem_interface is
    port (
        addr1,addr2 : in std_logic_vector (15 downto 0); -- addr1 is r/w, addr2 is r only
          wr_data : in std_logic_vector(15 downto 0);
          opcode : in std_logic_vector(6 downto 0);
          clk,rst : in std_logic;
          wr_en : in std_logic_vector(1 downto 0);
            r1_data,r2_data : out std_logic_vector(15 downto 0);
            err : out std_logic;
            disp_out : out std_logic_vector (15 downto 0); --for seven-seg-display
            in_port : in std_logic_vector(9 downto 0);
            out_port : out std_logic
    );
end component;

--IF/ID
component IF_ID is
    port (
        instr_in, pc_addr_in : in  std_logic_vector (15 downto 0);
        clk, rst, mem_stall : in  std_logic;
        pc_addr_out,op_pass : out std_logic_vector (15 downto 0);
        op_code: out std_logic_vector (6 downto 0);
        instr_format, reg1_addr, reg2_addr, ra_addr_out : out std_logic_vector (2 downto 0);
        mem_oper_out, wb_oper_out, m1_out : out std_logic
    );
end component;

--Register File
component register_file is
    port (
        rst : in std_logic; clk: in std_logic;
        --read signals
        rd_index1: in std_logic_vector(2 downto 0); 
        rd_index2: in std_logic_vector(2 downto 0); 
        rd_data1: out std_logic_vector(15 downto 0); 
        rd_data2: out std_logic_vector(15 downto 0);
        rd_vflag1: out std_logic;
        --write signals
        wr_index: in std_logic_vector(2 downto 0); 
        wr_data: in std_logic_vector(15 downto 0);
        wr_enable: in std_logic;
        v_flag: in std_logic
    );
end component;

--ID/EX
component ID_EX is 
    port (
        data_1, data_2, operand_3, pc_addr_in : in std_logic_vector (15 downto 0);
        opcode_in : in std_logic_vector (6 downto 0);
        instr_form_in, ra_addr_in, reg1_addr_in, reg2_addr_in : in std_logic_vector (2 downto 0);
        mem_oper_in, wb_oper_in, m1_in, v_flag_1, clk, rst, mem_stall : in std_logic;
        operand1, operand2, pc_addr_out, data_pass_out : out std_logic_vector (15 downto 0);
        opcode_out : out std_logic_vector (6 downto 0);
        alu_mode_out, instr_form_out, ra_addr_out, reg1_addr_out, reg2_addr_out : out std_logic_vector (2 downto 0);
        mem_oper_out, wb_oper_out, m1_out, v_flag_1_out : out std_logic
        );
end component;

--FWD_UNIT
component fwdunit is
    port(
        rst              : in STD_LOGIC;
        memwb_ra_addr    : in STD_LOGIC_VECTOR (2 downto 0);
        exmem_ra_addr    : in STD_LOGIC_VECTOR (2 downto 0);
        ifid_reg1_addr   : in STD_LOGIC_VECTOR (2 downto 0);
        ifid_reg2_addr   : in STD_LOGIC_VECTOR (2 downto 0);
        idex_reg1_addr   : in STD_LOGIC_VECTOR (2 downto 0);
        idex_reg2_addr   : in STD_LOGIC_VECTOR (2 downto 0);
        idex_ra_addr     : in STD_LOGIC_VECTOR (2 downto 0);
        idex_reg1_data   : in STD_LOGIC_VECTOR (15 downto 0);
        idex_reg2_data   : in STD_LOGIC_VECTOR (15 downto 0);
        idex_reg1_vflag  : in STD_LOGIC;
        idex_data_pass   : in STD_LOGIC_VECTOR (15 downto 0);
        idex_instr_form  : in STD_LOGIC_VECTOR (2 downto 0);
        idex_opcode_in   : in STD_LOGIC_VECTOR (6 downto 0);
        exmem_alu_result : in STD_LOGIC_VECTOR (15 downto 0);
        memwb_alu_result : in STD_LOGIC_VECTOR (15 downto 0);
        exmem_wb_oper    : in STD_LOGIC;
        memwb_wb_oper    : in STD_LOGIC;
        exmem_v_flag     : in STD_LOGIC;
        memwb_v_flag     : in STD_LOGIC;
        alu_operand1     : out STD_LOGIC_VECTOR (15 downto 0);
        alu_operand2     : out STD_LOGIC_VECTOR (15 downto 0);
        data_pass        : out STD_LOGIC_VECTOR (15 downto 0);
        v_flag_out       : out STD_LOGIC;
        stall_out        : out STD_LOGIC
    );
end component;

--ALU
component ALU is
    port (
        in1 : in std_logic_vector (15 downto 0);
        in2 : in std_logic_vector (15 downto 0);
        alu_mode : in std_logic_vector (2 downto 0);
        rst : in std_logic;
        result : out std_logic_vector (15 downto 0);
        z_flag : out std_logic;
        n_flag : out std_logic;
        v_flag : out std_logic
    );
end component;

--EX/MEM
component EX_MEM is
    port (
        alu_result, pc_addr_in, data_pass_in : in std_logic_vector (15 downto 0);
        opcode_in : in std_logic_vector (6 downto 0);
        instr_form_in, ra_addr_in : in std_logic_vector (2 downto 0);
        mem_oper_in, wb_oper_in, m1_in, clk, rst : in std_logic;
        alu_result_out, pc_addr_out, dest_data, src_data : out std_logic_vector (15 downto 0);
        opcode_out : out std_logic_vector (6 downto 0);
        instr_form_out, ra_addr_out : out std_logic_vector (2 downto 0);
        new_pc_addr_out: out std_logic_vector (15 downto 0);
        wb_oper_out : out std_logic;
        mem_oper_out : out std_logic_vector (1 downto 0);
        n_flag_in     : in std_logic; --Inputs from the status register, checked when branch instr reaches ex/mem
        z_flag_in    : in std_logic;
        v_flag_in      : in std_logic;
        v_flag_pass_in : in std_logic;
        br_flag_in   : in std_logic;
        br_trigger     : out std_logic;
        v_flag_pass_out: out std_logic
    );
end component;

--MEM/WB
component MEM_WB is 
    port (
        mem_data_in, alu_result_in, pc_addr_in : in std_logic_vector (15 downto 0);
        opcode_in : in std_logic_vector (6 downto 0);
        instr_format_in, ra_addr_in : in std_logic_vector (2 downto 0);
        wb_oper_in, clk, rst : in std_logic;
        v_flag_in     : in std_logic;
        wb_data_out   : out std_logic_vector (15 downto 0);
        ra_addr_out   : out std_logic_vector (2 downto 0);
        wb_oper_out   : out std_logic;
        v_flag_out    : out std_logic
    );
end component;

--STATUS REGISTER
component status_reg is
    port (clk, rst : in std_logic;
          n_flag_in : in std_logic;
          z_flag_in : in std_logic;
          v_flag_in : in std_logic;
          br_flag_in : in std_logic;
          clear_test_flags : in std_logic;
          n_flag_out : out std_logic;
          z_flag_out : out std_logic;
          v_flag_out : out std_logic;
          br_flag_out : out std_logic
    );
end component;

--DISPLAY CONTROLLER
component display_controller is
    port (clk, rst: in std_logic;
          hex3, hex2, hex1, hex0: in std_logic_vector(3 downto 0);
          an: out std_logic_vector(3 downto 0);
          sseg: out std_logic_vector(6 downto 0)   
          );
end component;
-- Constants
constant instr_mem_size : integer := 2; -- each instr is 2 bytes

--GLOBAL
signal clk_sig   : std_logic;
signal rst : std_logic;
signal rst_sig   : std_logic := '0';
signal stall_sig : std_logic := '0';
signal rl_flag :std_logic := '0';
signal re_flag :std_logic := '0';

--INSTRUCTION FETCH
signal instr_mem_output : std_logic_vector (15 downto 0) := (others => '0');
signal ifid_pc_addr_out : std_logic_vector (15 downto 0):= (others => '0');
signal ifid_op_pass_out : std_logic_vector (15 downto 0):= (others => '0');
signal ifid_opcode_out : std_logic_vector (6 downto 0):= (others => '0');
signal ifid_instr_format_out : std_logic_vector (2 downto 0):= (others => '0');
signal ifid_reg1_addr_out : std_logic_vector (2 downto 0):= (others => '0');
signal ifid_reg2_addr_out : std_logic_vector (2 downto 0):= (others => '0');
signal if_id_ra_addr_out  : std_logic_vector (2 downto 0):= (others => '0');
signal ifid_mem_oper_out : std_logic := '0';
signal ifid_wb_oper_out : std_logic := '0';
signal ifid_m1_out : std_logic := '0';

--INSTRUCTION DECODE
signal regfile_reg1_data_out : std_logic_vector (15 downto 0);
signal regfile_reg2_data_out : std_logic_vector (15 downto 0);
signal regfile_reg1_v_flag : std_logic;
signal idex_reg1_data_out : std_logic_vector (15 downto 0):= (others => '0');
signal idex_reg2_data_out : std_logic_vector (15 downto 0):= (others => '0');
signal idex_opcode_out : std_logic_vector (6 downto 0):= (others => '0');
signal idex_alu_mode_out : std_logic_vector (2 downto 0):= (others => '0');
signal idex_instr_form_out : std_logic_vector (2 downto 0):= (others => '0');
signal idex_pc_addr_out : std_logic_vector (15 downto 0):= (others => '0');
signal idex_data_pass_out : std_logic_vector (15 downto 0):= (others => '0');
signal idex_ra_addr_out : std_logic_vector (2 downto 0):= (others => '0');
signal idex_r1_addr_out : std_logic_vector (2 downto 0):= (others => '0');
signal idex_r2_addr_out : std_logic_vector (2 downto 0):= (others => '0');
signal idex_mem_oper_out : std_logic;
signal idex_wb_oper_out : std_logic;
signal idex_m1_out : std_logic := '0';
signal idex_vflag_out : std_logic := '0';

signal fwd_unit_operand1_out : std_logic_vector (15 downto 0):= (others => '0');
signal fwd_unit_operand2_out : std_logic_vector (15 downto 0):= (others => '0');
signal fwd_unit_data_pass_out : std_logic_vector (15 downto 0):= (others => '0');
signal fwd_unit_vflag_out : std_logic:= '0';

--EXECUTE
signal alu_result_out : std_logic_vector (15 downto 0):= (others => '0');
signal alu_z_flag_out : std_logic;
signal alu_n_flag_out : std_logic;
signal alu_v_flag_out : std_logic;
signal exmem_alu_result_out : std_logic_vector (15 downto 0):= (others => '0');
signal exmem_pc_addr_out : std_logic_vector (15 downto 0):= (others => '0');
signal exmem_dest_data_out : std_logic_vector (15 downto 0):= (others => '0');
signal exmem_src_data_out : std_logic_vector (15 downto 0):= (others => '0');
signal exmem_opcode_out : std_logic_vector (6 downto 0):= (others => '0');
signal exmem_instr_form_out : std_logic_vector (2 downto 0):= (others => '0');
signal exmem_ra_addr_out : std_logic_vector (2 downto 0):= (others => '0');
signal exmem_mem_oper_out : std_logic_vector (1 downto 0):= (others => '0');
signal exmem_wb_oper_out : std_logic;
signal exmem_vflag_out : std_logic:= '0';

--MEMORY/WB
signal data_mem_output : std_logic_vector (15 downto 0):= (others => '0');
signal memwb_data_out : std_logic_vector (15 downto 0):= (others => '0');
signal memwb_ra_addr_out : std_logic_vector (2 downto 0):= (others => '0');
signal memwb_wb_oper_out : std_logic:= '0';
signal memwb_vflag_out : std_logic:= '0';

--BRANCHING
signal exmem_br_addr_out : std_logic_vector (15 downto 0) := (others => '0');
signal exmem_br_trig_out : std_logic := '0';

--PC behaviour
signal pc_addr : std_logic_vector(15 downto 0):= (others => '0');
signal pc_next_addr : std_logic_vector(15 downto 0):= (others => '0');

--STATUS REGISTER
signal stat_reg_n_out : std_logic;
signal stat_reg_z_out : std_logic;
signal stat_reg_v_out : std_logic;
signal stat_reg_br_out : std_logic;
signal stat_reg_clr_flag_in : std_logic;

--DISPLAY
signal sw_sig : std_logic_vector(1 downto 0) := (others => '0');
signal disp_out : std_logic_vector(15 downto 0) := (others => '0');

begin
-- Component port mappings

--PC
pc0 : pc port map (
    clk => clk,
    rst => rst_sig,
    pc_in => pc_next_addr,
    pc_out => pc_addr
);

--Mem Module
mem0 : mem_interface port map (
    clk => clk,
    rst => rst_sig,
    err => open,
    
    --INSTRUCTION MEMORY
    addr2 => pc_addr,
    r2_data => instr_mem_output,

    --DATA MEMORY
    addr1 => exmem_dest_data_out,
    wr_data => exmem_src_data_out,
    wr_en => exmem_mem_oper_out,
    r1_data => data_mem_output,
    
    --INPUT AND OUTPUT PORTS
    in_port => in_port,
    out_port => out_port,
    opcode => exmem_opcode_out,
    disp_out => disp_out
);

--IF/ID
ifid0: if_id port map(
    clk => clk,
    rst => rst_sig,
    mem_stall => stall_sig,
    
    instr_in => instr_mem_output,
    pc_addr_in => pc_addr,
    
    pc_addr_out => ifid_pc_addr_out,
    op_pass => ifid_op_pass_out,
    op_code => ifid_opcode_out,
    instr_format => ifid_instr_format_out,
    reg1_addr => ifid_reg1_addr_out,
    reg2_addr => ifid_reg2_addr_out,
    mem_oper_out => ifid_mem_oper_out,
    wb_oper_out => ifid_wb_oper_out,
    m1_out => ifid_m1_out,
    ra_addr_out => if_id_ra_addr_out
);

--Reg File
rf0: register_file port map (
    clk => clk,
    rst => rst,
    
    --READ
    rd_index1 => ifid_reg1_addr_out,
    rd_index2 => ifid_reg2_addr_out,
    rd_data1 => regfile_reg1_data_out,
    rd_data2 => regfile_reg2_data_out,
    rd_vflag1 => regfile_reg1_v_flag,
    
    --WRITE
    wr_index => memwb_ra_addr_out,
    wr_data => memwb_data_out,
    wr_enable => memwb_wb_oper_out,
    v_flag => memwb_vflag_out
);

--ID/EX
idex0 : id_ex port map (
    clk => clk,
    rst => rst_sig,
    mem_stall => stall_sig,
    
    data_1 => regfile_reg1_data_out,
    data_2 => regfile_reg2_data_out,
    v_flag_1 => regfile_reg1_v_flag,
    operand_3 => ifid_op_pass_out,
    opcode_in => ifid_opcode_out,
    instr_form_in => ifid_instr_format_out,
    ra_addr_in => if_id_ra_addr_out,
    reg1_addr_in => ifid_reg1_addr_out,
    reg2_addr_in => ifid_reg2_addr_out,
    pc_addr_in => ifid_pc_addr_out,
    mem_oper_in => ifid_mem_oper_out,
    wb_oper_in => ifid_wb_oper_out,
    m1_in => ifid_m1_out,
    operand1 => idex_reg1_data_out,
    operand2 => idex_reg2_data_out,

    opcode_out => idex_opcode_out,
    alu_mode_out => idex_alu_mode_out,
    instr_form_out => idex_instr_form_out,
    pc_addr_out => idex_pc_addr_out,
    data_pass_out => idex_data_pass_out,
    ra_addr_out => idex_ra_addr_out,
    reg1_addr_out => idex_r1_addr_out,
    reg2_addr_out => idex_r2_addr_out,
    mem_oper_out => idex_mem_oper_out,
    wb_oper_out => idex_wb_oper_out,
    m1_out => idex_m1_out,
    v_flag_1_out => idex_vflag_out
);

--FWD_UNIT
fu0: fwdunit port map (
    rst => rst_sig,
    ifid_reg1_addr => ifid_reg1_addr_out,
    ifid_reg2_addr => ifid_reg2_addr_out,
    idex_ra_addr => idex_ra_addr_out,
    idex_reg1_data => idex_reg1_data_out,
    idex_reg2_data => idex_reg2_data_out,
    idex_reg1_vflag => idex_vflag_out,
    idex_data_pass => idex_data_pass_out,
    idex_reg1_addr => idex_r1_addr_out,
    idex_reg2_addr => idex_r2_addr_out,
    idex_instr_form => idex_instr_form_out,
    idex_opcode_in => idex_opcode_out,
    exmem_alu_result => exmem_alu_result_out,
    memwb_alu_result => memwb_data_out,
    exmem_wb_oper => exmem_wb_oper_out,
    memwb_wb_oper => memwb_wb_oper_out,
    exmem_v_flag => exmem_vflag_out,
    memwb_v_flag => memwb_vflag_out,
    exmem_ra_addr => exmem_ra_addr_out,
    memwb_ra_addr => memwb_ra_addr_out,
    
    alu_operand1 => fwd_unit_operand1_out,
    alu_operand2 => fwd_unit_operand2_out,
    data_pass => fwd_unit_data_pass_out,
    v_flag_out => fwd_unit_vflag_out,
    stall_out => stall_sig
);


--ALU
alu0: alu port map (
    rst => rst_sig,
    in1 => fwd_unit_operand1_out,
    in2 => fwd_unit_operand2_out,
    alu_mode => idex_alu_mode_out,
    result => alu_result_out,
    z_flag => alu_z_flag_out,
    n_flag => alu_n_flag_out,
    v_flag => alu_v_flag_out
);

--EX/MEM
exmem0: ex_mem port map (
    clk => clk,
    rst => rst,

    alu_result => alu_result_out,
    instr_form_in => idex_instr_form_out,
    opcode_in => idex_opcode_out,
    pc_addr_in => idex_pc_addr_out,
    data_pass_in => fwd_unit_data_pass_out,
    ra_addr_in => idex_ra_addr_out,
    mem_oper_in => idex_mem_oper_out,
    wb_oper_in => idex_wb_oper_out,
    m1_in => idex_m1_out,
    n_flag_in => stat_reg_n_out,
    z_flag_in => stat_reg_z_out,
    v_flag_in => stat_reg_v_out,
    v_flag_pass_in => alu_v_flag_out,
    br_flag_in => stat_reg_br_out,
    
    alu_result_out => exmem_alu_result_out,
    pc_addr_out => exmem_pc_addr_out,
    dest_data => exmem_dest_data_out,
    src_data => exmem_src_data_out,
    opcode_out => exmem_opcode_out,
    instr_form_out => exmem_instr_form_out,
    ra_addr_out => exmem_ra_addr_out,
    mem_oper_out => exmem_mem_oper_out,
    wb_oper_out => exmem_wb_oper_out,
    v_flag_pass_out => exmem_vflag_out,
    br_trigger => exmem_br_trig_out,
    new_pc_addr_out => exmem_br_addr_out
);

--MEM/WB
memwb0: mem_wb port map (
    clk => clk,
    rst => rst,

    mem_data_in => data_mem_output,
    alu_result_in => exmem_alu_result_out,
    instr_format_in => exmem_instr_form_out,
    pc_addr_in => exmem_pc_addr_out,
    opcode_in => exmem_opcode_out,
    ra_addr_in => exmem_ra_addr_out,
    wb_oper_in => exmem_wb_oper_out,
    v_flag_in => exmem_vflag_out,
    
    wb_data_out => memwb_data_out,
    ra_addr_out => memwb_ra_addr_out,
    wb_oper_out => memwb_wb_oper_out,
    v_flag_out => memwb_vflag_out
    
);

--STATUS REGISTER
sr0: status_reg port map (
     clk => clk,
     rst => rst,
     n_flag_in => alu_n_flag_out,
     z_flag_in => alu_z_flag_out,
     v_flag_in => fwd_unit_vflag_out,
     br_flag_in => exmem_br_trig_out,
     clear_test_flags => stat_reg_clr_flag_in,
     n_flag_out => stat_reg_n_out,
     z_flag_out => stat_reg_z_out,
     v_flag_out => stat_reg_v_out,
     br_flag_out => stat_reg_br_out
);

--DISPLAY
dc0: display_controller port map (
    clk => clk,
    rst => rst,
    hex3 => disp_out(15 downto 12),
    hex2 => disp_out(11 downto 8),
    hex1 => disp_out(7 downto 4),
    hex0 => disp_out(3 downto 0),
    an => an_out,
    sseg => sseg_out
);

           

--Combinational logic
    -- Detected branch, 
    -- if BR.SUB, store the PC_address in r7 and use new pc addr from R[ra]
    -- r7 <= exmem_pc_addr_out + instr_mem_size
    -- (store incremented address)
    
    rl_flag <= sw_in(0);
    re_flag <= sw_in(1);

    rst <= (sw_in(0) or sw_in(1));
    
    pc_next_addr <= (others => '0') when rst_sig = '1' else 
		    exmem_br_addr_out when exmem_br_trig_out = '1' else
		    pc_addr when stall_sig = '1' else
		    X"0002" when sw_in(0) = '1' else --Load
		    X"0000" when sw_in(1) = '1' else --Exe
            std_logic_vector(unsigned(pc_addr) + instr_mem_size);
    
    --set clear on succesful branch
    stat_reg_clr_flag_in <= '1' when stat_reg_br_out = '1' else '0';
    
    rst_sig <= '1' when exmem_br_trig_out = '1' else -- reset if/id and id/ex when branching
               rst; -- follow processor reset otherwise
                

   
    --STALL BEHAVIOUR

end behavioral;
