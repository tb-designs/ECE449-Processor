
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity incrementor is


end incrementor;