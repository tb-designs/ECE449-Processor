library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity MEM_WB is 
  port();

end MEM_WB;

architecture Behavioral of MEM_WB is


  end Behavioral;