library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity EX_MEM is 
  port();

end EX_MEM;

architecture Behavioral of EX_MEM is


  end Behavioral;